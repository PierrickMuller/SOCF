-----------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- File         : axi4lite_slave.vhd
-- Author       : E. Messerli    27.07.2017
-- Description  : slave interface AXI  (without burst)
-- used for     : SOCF lab
--| Modifications |-----------------------------------------------------------
-- Ver  Date       Auteur  Description
-- 1.0  26.03.2019  EMI    Adaptation du chablon pour les etudiants  
--
------------------------------------------------------------------------------
-- Pas utiliser les deux bits de poids faible


library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

entity axi4lite_slave is
    generic (
        -- Users to add parameters here

        -- User parameters ends

        -- Width of S_AXI data bus
        AXI_DATA_WIDTH  : integer   := 32;  -- 32 or 64 bits
        -- Width of S_AXI address bus
        AXI_ADDR_WIDTH  : integer   := 12
    );
    port (
        axi_clk_i       : in  std_logic;
        axi_reset_i     : in  std_logic;
        -- AXI4-Lite 
        axi_awaddr_i    : in  std_logic_vector(AXI_ADDR_WIDTH-1 downto 0);
        axi_awprot_i    : in  std_logic_vector( 2 downto 0); -- Pas utilisés
        axi_awvalid_i   : in  std_logic;
        axi_awready_o   : out std_logic;
        axi_wdata_i     : in  std_logic_vector(AXI_DATA_WIDTH-1 downto 0);
        axi_wstrb_i     : in std_logic_vector((AXI_DATA_WIDTH/8)-1 downto 0); -- A gérer aussi 
        axi_wvalid_i    : in  std_logic;
        axi_wready_o    : out std_logic;
        axi_bresp_o     : out std_logic_vector(1 downto 0);
        axi_bvalid_o    : out std_logic;
        axi_bready_i    : in  std_logic;
        axi_araddr_i    : in  std_logic_vector(AXI_ADDR_WIDTH-1 downto 0);
        axi_arprot_i    : in  std_logic_vector( 2 downto 0); -- Pas utilisés
        axi_arvalid_i   : in  std_logic;
        axi_arready_o   : out std_logic;
        axi_rdata_o     : out std_logic_vector(AXI_DATA_WIDTH-1 downto 0);
        axi_rresp_o     : out std_logic_vector(1 downto 0);
        axi_rvalid_o    : out std_logic;
        axi_rready_i    : in  std_logic
        -- User input-output
        
        
    );
end entity axi4lite_slave;

architecture rtl of axi4lite_slave is

    signal reset_s : std_logic;

    -- local parameter for addressing 32 bit / 64 bits, cst: AXI_DATA_WIDTH
    -- ADDR_LSB is used for addressing word 32/64 bits registers/memories
    -- ADDR_LSB = 2 for 32 bits (n-1 downto 2)
    -- ADDR_LSB = 3 for 64 bits (n-1 downto 3)
    constant ADDR_LSB  : integer := (AXI_DATA_WIDTH/32)+ 1;
    
    --signal for the AXI slave
    --intern signal for output
    signal axi_awready_s       : std_logic;
    signal axi_arready_s       : std_logic;

     --intern signal for the axi interface
    signal axi_waddr_mem_s     : std_logic_vector(AXI_ADDR_WIDTH-1 downto ADDR_LSB);
    signal axi_araddr_mem_s    : std_logic_vector(AXI_ADDR_WIDTH-1 downto ADDR_LSB);
    
     --intern signal for adress decoding
    signal local_address_write_s <=    : integer;
    signal local_address_read_s <=	  : integer;
	signal const_register_address_valid_write_s : std_logic;
	signal test_register_address_valid_write_s : std_logic;
	signal leds_register_address_valid_write_s : std_logic;
	signal hex03_register_address_valid_write_s : std_logic;
	signal hex45_register_address_valid_write_s : std_logic;
	signal switch_register_address_valid_write_s : std_logic;
	signal keys_register_address_valid_write_s : std_logic;
	signal const_register_address_valid_read_s : std_logic;
	signal test_register_address_valid_read_s : std_logic;
	signal leds_register_address_valid_read_s : std_logic;
	signal hex03_register_address_valid_read_s : std_logic;
	signal hex45_register_address_valid_read_s : std_logic;
	signal switch_register_address_valid_read_s : std_logic;
	signal keys_register_address_valid_read_s : std_logic;
begin

    reset_s  <= axi_reset_i;

-----------------------------------------------------------
-- address decoding

-- On récupére l'offset dans l'adresse. On utilise pas les deux bits de poid faible 
local_address_write_s <= to_integer(unsigned(axi_waddr_mem_s(AXI_ADDR_WIDTH - 1 downto 0)));
local_address_read_s <= to_integer(unsigned(axi_araddr_mem_s(AXI_ADDR_WIDTH - 1 downto 0)));

address_range_analysis : process (local_address_write_s, local_address_read_s)
begin
	-- write valid
	const_register_address_valid_write_s <= '0';
	test_register_address_valid_write_s <= '0';
	leds_register_address_valid_write_s <= '0';
	hex03_register_address_valid_write_s <= '0';
	hex45_register_address_valid_write_s <= '0';
	switch_register_address_valid_write_s <= '0';
	keys_register_address_valid_write_s <= '0';
	
	-- read valid 
	const_register_address_valid_read_s <= '0';
	test_register_address_valid_read_s <= '0';
	leds_register_address_valid_read_s <= '0';
	hex03_register_address_valid_read_s <= '0';
	hex45_register_address_valid_read_s <= '0';
	switch_register_address_valid_read_s <= '0';
	keys_register_address_valid_read_s <= '0';	
	
	case (local_address_write_s) is
		when 0 => const_register_address_valid_write_s <= '1';
		when 1 => test_register_address_valid_write_s <= '1';
		when 2 => leds_register_address_valid_write_s <= '1'; 
		when 3 => hex03_register_address_valid_write_s <= '1';
		when 4 => hex45_register_address_valid_write_s <= '1';
		when 5 => switch_register_address_valid_write_s <= '1';
		when 6 => keys_register_address_valid_write_s <= '1';
		when others => NULL;
	end case;
	
	case (local_address_read_s) is
		when 0 => const_register_address_valid_read_s <= '1';
		when 1 => test_register_address_valid_read_s <= '1';
		when 2 => leds_register_address_valid_read_s <= '1'; 
		when 3 => hex03_register_address_valid_read_s <= '1';
		when 4 => hex45_register_address_valid_read_s <= '1';
		when 5 => switch_register_address_valid_read_s <= '1';
		when 6 => keys_register_address_valid_read_s <= '1';
		when others => NULL;
	end case;
end process;

-----------------------------------------------------------
-- Write address channel

    process (reset_s, axi_clk_i)
    begin
        if reset_s = '1' then
            axi_awready_s <= '0';
            axi_waddr_mem_s <= (others => '0');
        elsif rising_edge(axi_clk_i) then
            if (axi_awready_s = '0' and axi_awvalid_i = '1')  then --and axi_wvalid_i = '1') then  modif EMI 10juil2018
                -- slave is ready to accept write address when
                -- there is a valid write address
                axi_awready_s <= '1';
                -- Write Address memorizing
                axi_waddr_mem_s <= axi_awaddr_i(AXI_ADDR_WIDTH-1 downto ADDR_LSB);
            else
                axi_awready_s <= '0';
            end if;
        end if;
    end process;
    axi_awready_o <= axi_awready_s;


-----------------------------------------------------------
-- Write data channel

    -- Implement axi_wready generation
    process (reset_s, clk_i)
    begin
        if reset_s = '1' then
            axi_waddr_done_s <= '0'; 
            axi_wready_s    <= '0';
        elsif rising_edge(clk_i) then

        
          --to be completed
           
        
        
        end if;
    end process;
    
    axi_wready_o <= axi_wready_s;


    --condition to write data
    axi_data_wren_s <=  --to be completed....     ;
    
    
    process (reset_s, clk_i)
        --number address to access 32 or 64 bits data
        variable int_waddr_v : natural;
    begin
        if reset_s = '1' then
            
          --to be completed
            
            
        elsif rising_edge(clk_i) then

            if axi_data_wren_s = '1' then
                int_waddr_v   := to_integer(unsigned(axi_waddr_mem_s));
                case int_waddr_v is
                    when 0   => .....
                    
                    when 1   => .....
                    
                    
                    --to be completed


                    when others => null;
                end case;
            end if;
        end if;
    end process;
                    

-----------------------------------------------------------
-- Write response channel


    --to be completed


    

-----------------------------------------------------------
-- Read address channel

    process (reset_s, axi_clk_i)
    begin
        if reset_s = '1' then
           axi_arready_s    <= '0';
           axi_araddr_mem_s <= (others => '1');
        elsif rising_edge(axi_clk_i) then
            if axi_arready_s = '0' and axi_arvalid_i = '1' then
                -- indicates that the slave has acceped the valid read address
                axi_arready_s    <= '1';
                -- Read Address memorizing
                axi_araddr_mem_s <= axi_araddr_i(AXI_ADDR_WIDTH-1 downto ADDR_LSB);
            else
                axi_arready_s    <= '0';
            end if;
        end if;
    end process;
    axi_arready_o <= axi_arready_s;

-----------------------------------------------------------
-- Read data channel

    --to be completed



end rtl;
